module main

println('vlang is able to write like this (no fn main()).')
